module hello_world();

initial begin
 $display("\n\t Hello world! \n");
end

endmodule